module Lab3bUnMinimized(
input a,
input b,
input c,
output out
);
bc
abc
endmodule
