module Lab3bMinimized(
input a,
input b,
input c,
output out
);
bc
endmodule
